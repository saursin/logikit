`define UNUSED_VAR(x) always @(x) begin end